--Jonathan Cruz
--University of Florida

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants.all;

entity round is
    port(
        x	: in std_logic_vector(WORD_SIZE-1 downto 0); --most significant word of input
        y	: in std_logic_vector(WORD_SIZE-1 downto 0); -- least signficant word of input
	round_key : in std_logic_vector(WORD_SIZE-1 downto 0); 
	round_out : out std_logic_vector(BLOCK_SIZE-1 downto 0)
    );

end round;

architecture BHV of round is


begin
    process(x,y,round_key)
	----------- your variables here -----------
	
    begin
	----------- your code here -----------

	
    end process;
end BHV;
